module control
(
	input logic [5:0] opcode,
	input logic [5:0] func,
	input logic zero,
	output logic [12:0] control
);

endmodule